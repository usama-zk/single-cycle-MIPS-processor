`timescale 1ns / 1ps
module Regfile(clk,RegWrite,rs,rt,rd,rs_out,rt_out,rd_in);
input clk,RegWrite;
input [4:0] rs,rt,rd;
output reg [31:0] rs_out,rt_out;
input [31:0] rd_in;
reg [31:0] mem[31:0];
initial
begin
mem[0]=32'd5;
mem[1]=32'd10;
mem[2]=32'd20;
mem[3]=32'd25;
mem[4]=32'd30;
mem[5]=32'd35;
mem[6]=32'd40;
mem[7]=32'd45;
mem[8]=32'd50;
mem[9]=32'd55;
mem[10]=32'd60;
mem[11]=32'd65;
mem[12]=32'd70;
mem[13]=32'd75;
mem[14]=32'd80;
mem[15]=32'd85;
mem[16]=32'd90;
mem[17]=32'd95;
mem[18]=32'd100;
mem[19]=32'd105;
mem[20]=32'd110;
mem[21]=32'd115;
mem[22]=32'd120;
mem[23]=32'd125;
mem[24]=32'd130;
mem[25]=32'd135;
mem[26]=32'd140;
mem[27]=32'd145;
mem[28]=32'd150;
mem[29]=32'd155;
mem[30]=32'd160;
mem[31]=32'd165;
end


always @(*)
begin
case(rs)
32'd0:rs_out<=mem[0];
32'd1:rs_out<=mem[1];
32'd2:rs_out<=mem[2];
32'd3:rs_out<=mem[3];
32'd4:rs_out<=mem[4];
32'd5:rs_out<=mem[5];
32'd6:rs_out<=mem[6];
32'd7:rs_out<=mem[7];
32'd8:rs_out<=mem[8];
32'd9:rs_out<=mem[9];
32'd10:rs_out<=mem[10];
32'd11:rs_out<=mem[11];
32'd12:rs_out<=mem[12];
32'd13:rs_out<=mem[13];
32'd14:rs_out<=mem[14];
32'd15:rs_out<=mem[15];
32'd16:rs_out<=mem[16];
32'd17:rs_out<=mem[17];
32'd18:rs_out<=mem[18];
32'd19:rs_out<=mem[19];
32'd20:rs_out<=mem[20];
32'd21:rs_out<=mem[21];
32'd22:rs_out<=mem[22];
32'd23:rs_out<=mem[23];
32'd24:rs_out<=mem[24];
32'd25:rs_out<=mem[25];
32'd26:rs_out<=mem[26];
32'd27:rs_out<=mem[27];
32'd28:rs_out<=mem[28];
32'd29:rs_out<=mem[29];
32'd30:rs_out<=mem[30];
32'd31:rs_out<=mem[31];
endcase
case(rt)
32'd0:rt_out<=mem[0];
32'd1:rt_out<=mem[1];
32'd2:rt_out<=mem[2];
32'd3:rt_out<=mem[3];
32'd4:rt_out<=mem[4];
32'd5:rt_out<=mem[5];
32'd6:rt_out<=mem[6];
32'd7:rt_out<=mem[7];
32'd8:rt_out<=mem[8];
32'd9:rt_out<=mem[9];
32'd10:rt_out<=mem[10];
32'd11:rt_out<=mem[11];
32'd12:rt_out<=mem[12];
32'd13:rt_out<=mem[13];
32'd14:rt_out<=mem[14];
32'd15:rt_out<=mem[15];
32'd16:rt_out<=mem[16];
32'd17:rt_out<=mem[17];
32'd18:rt_out<=mem[18];
32'd19:rt_out<=mem[19];
32'd20:rt_out<=mem[20];
32'd21:rt_out<=mem[21];
32'd22:rt_out<=mem[22];
32'd23:rt_out<=mem[23];
32'd24:rt_out<=mem[24];
32'd25:rt_out<=mem[25];
32'd26:rt_out<=mem[26];
32'd27:rt_out<=mem[27];
32'd28:rt_out<=mem[28];
32'd29:rt_out<=mem[29];
32'd30:rt_out<=mem[30];
32'd31:rt_out<=mem[31];
endcase

if(RegWrite)
case(rd)
32'd0:mem[0]<=rd_in;
32'd1:mem[1]<=rd_in;
32'd2:mem[2]<=rd_in;
32'd3:mem[3]<=rd_in;
32'd4:mem[4]<=rd_in;
32'd5:mem[5]<=rd_in;
32'd6:mem[6]<=rd_in;
32'd7:mem[7]<=rd_in;
32'd8:mem[8]<=rd_in;
32'd9:mem[9]<=rd_in;
32'd10:mem[10]<=rd_in;
32'd11:mem[11]<=rd_in;
32'd12:mem[12]<=rd_in;
32'd13:mem[13]<=rd_in;
32'd14:mem[14]<=rd_in;
32'd15:mem[15]<=rd_in;
32'd16:mem[16]<=rd_in;
32'd17:mem[17]<=rd_in;
32'd18:mem[18]<=rd_in;
32'd19:mem[19]<=rd_in;
32'd20:mem[20]<=rd_in;
32'd21:mem[21]<=rd_in;
32'd22:mem[22]<=rd_in;
32'd23:mem[23]<=rd_in;
32'd24:mem[24]<=rd_in;
32'd25:mem[25]<=rd_in;
32'd26:mem[26]<=rd_in;
32'd27:mem[27]<=rd_in;
32'd28:mem[28]<=rd_in;
32'd29:mem[29]<=rd_in;
32'd30:mem[30]<=rd_in;
32'd31:mem[31]<=rd_in;
endcase
end
endmodule
