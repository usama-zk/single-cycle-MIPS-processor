`timescale 1ns / 1ps
module Jump_Ext(J_in,J_out);
input [25:0] J_in;
output reg [31:0] J_out;


endmodule
